** sch_path: /foss/designs/ADT_Designs/cs_stage.sch
**.subckt cs_stage Vout
*.opin Vout
V1 vdd GND 1.8
R1 vdd Vout 100k m=1
I0 vdd net1 10u
XM4 net1 net1 GND GND sg13_hv_nmos w=2.8u l=2u ng=1 m=1
R7 net2 net1 1 ac=1e12 m=1
R8 net3 net2 1e12 ac=1 m=1
V2 net3 GND DC 0 AC 1
XM1 Vout net2 GND GND sg13_lv_nmos w=1.0u l=0.45u ng=1 m=1
**** begin user architecture code



.lib cornerMOSlv.lib mos_tt
.lib cornerMOShv.lib mos_tt
.lib cornerHBT.lib hbt_typ
.lib cornerRES.lib res_typ





.control
save all
op
write cs_stage.raw
ac dec 10 1 10g
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
